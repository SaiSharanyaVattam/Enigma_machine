`timescale 1ns / 1ps

module USB_Receiver(
    input clk,
    input kclk,
    input kdata,
    output reg [15:0] keycode=0,
    output reg oflag,
    output myflag
    );

    wire kclkf, kdataf;
    reg [7:0]datacur=0;
    reg [7:0]dataprev=0;
    reg [3:0]cnt=0;
    reg flag=0;
    //reg temp = 0;
//    initial begin
//        myflag = 0;
//    end


    debouncer #(
        .COUNT_MAX(19),
        .COUNT_WIDTH(5)
    ) db_clk(
        .clk(clk),
        .I(kclk),
        .O(kclkf)
    );
    debouncer #(
       .COUNT_MAX(19),
       .COUNT_WIDTH(5)
    ) db_data(
        .clk(clk),
        .I(kdata),
        .O(kdataf)
    );
    assign myflag = kdataf;
    always@(negedge(kclkf))begin
        case(cnt)
        0:;//Start bit
        1:datacur[0]<=kdataf;
        2:datacur[1]<=kdataf;
        3:datacur[2]<=kdataf;
        4:datacur[3]<=kdataf;
        5:datacur[4]<=kdataf;
        6:datacur[5]<=kdataf;
        7:datacur[6]<=kdataf;
        8:datacur[7]<=kdataf;
        9:flag<=1'b1;
        10:flag<=1'b0;
    
        endcase
            if(cnt<=9) cnt<=cnt+1;
            else if(cnt==10) cnt<=0;
    end
    
    reg pflag;
    always@(posedge clk) begin
        if (flag == 1'b1 && pflag == 1'b0) begin
            keycode <= {dataprev, datacur};
            oflag <= 1'b1;
            dataprev <= datacur;
            //temp <= 1;
            //myflag <= 1'b1;
        end else
            oflag <= 'b0;
        pflag <= flag;
    end

endmodule
